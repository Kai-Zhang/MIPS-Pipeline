module ControlHazard(
output reg Keep,
output reg Reset
);
initial 
begin 
Keep=0;
Reset=0;
end 
endmodule
