library verilog;
use verilog.vl_types.all;
entity ID_Ex is
    port(
        clk             : in     vl_logic;
        Reset           : in     vl_logic;
        Rs_in           : in     vl_logic_vector(4 downto 0);
        Rt_in           : in     vl_logic_vector(4 downto 0);
        Rd_in           : in     vl_logic_vector(4 downto 0);
        Rs_out_in       : in     vl_logic_vector(31 downto 0);
        Rt_out_in       : in     vl_logic_vector(31 downto 0);
        offset_in       : in     vl_logic_vector(31 downto 0);
        RegDst_in       : in     vl_logic;
        Shift_amountSrc_in: in     vl_logic;
        Jump_in         : in     vl_logic;
        ALUShift_Sel_in : in     vl_logic;
        RegDt0_in       : in     vl_logic;
        ALU_op_in       : in     vl_logic_vector(3 downto 0);
        Shift_op_in     : in     vl_logic_vector(1 downto 0);
        ALUSrcB_in      : in     vl_logic_vector(1 downto 0);
        Condition_in    : in     vl_logic_vector(2 downto 0);
        LoadType_in     : in     vl_logic_vector(1 downto 0);
        LoadByte_in     : in     vl_logic_vector(1 downto 0);
        RegWr_in        : in     vl_logic;
        MemWr_in        : in     vl_logic;
        MemtoReg_in     : in     vl_logic;
        PC_in           : in     vl_logic_vector(31 downto 0);
        Target_in       : in     vl_logic_vector(25 downto 0);
        Shamt_in        : in     vl_logic_vector(4 downto 0);
        Rs_out          : out    vl_logic_vector(4 downto 0);
        Rt_out          : out    vl_logic_vector(4 downto 0);
        Rd_out          : out    vl_logic_vector(4 downto 0);
        Rs_out_out      : out    vl_logic_vector(31 downto 0);
        Rt_out_out      : out    vl_logic_vector(31 downto 0);
        offset_out      : out    vl_logic_vector(31 downto 0);
        RegDst_out      : out    vl_logic;
        Shift_amountSrc_out: out    vl_logic;
        Jump_out        : out    vl_logic;
        ALUShift_Sel_out: out    vl_logic;
        RegDt0_out      : out    vl_logic;
        ALU_op_out      : out    vl_logic_vector(3 downto 0);
        Shift_op_out    : out    vl_logic_vector(1 downto 0);
        ALUSrcB_out     : out    vl_logic_vector(1 downto 0);
        Condition_out   : out    vl_logic_vector(2 downto 0);
        LoadType_out    : out    vl_logic_vector(1 downto 0);
        LoadByte_out    : out    vl_logic_vector(1 downto 0);
        RegWr_out       : out    vl_logic;
        MemWr_out       : out    vl_logic;
        MemtoReg_out    : out    vl_logic;
        PC_out          : out    vl_logic_vector(31 downto 0);
        Target_Out      : out    vl_logic_vector(25 downto 0);
        Shamt_out       : out    vl_logic_vector(4 downto 0)
    );
end ID_Ex;
